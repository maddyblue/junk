* potentiostat
.options  tnom=27
.temp 27

* OPA827 - operational amplifier SPICE MODEL
*
* Amplifier classification: Low-noise, high-precision, JFET-input, operational amplifier
*
* Model Definition by T E Kuehl - Texas Instruments Inc.
*
* Rev. A - 26 September 2008, by W.K. SANDS
*
*     This macromodel has been optimized to model the AC, DC, noise, and transient response performance within
*     the device data sheet specified limits. Correct operation of this macromodel has been verified on
*     MicroSim P-Spice ver. 8.0, DesignSoft TINA, and on PENZAR Development TopSPICE ver. 6.82d. For help
*     with other analog simulation software, please consult your software supplier.
*
* Copyright 2008 by Texas Instruments Corporation
*
* BEGIN MODEL OPA827
* PINOUT ORDER +IN -IN +V -V OUT
* PINOUT ORDER  3   2   7  4  6
.SUBCKT OPA827 3 2 7 4 6
* BEGIN MODEL FEATURES
* OPEN LOOP GAIN AND PHASE, INPUT OFFSET VOLTAGE W TEMPCO,
* INPUT VOLTAGE NOISE WITH 1/F, INPUT CURRENT NOISE, INPUT
* BIAS CURRENT W TEMPERATURE EFFECTS, INPUT CAPACITANCE,
* INPUT COMMON MODE VOLTAGE RANGE, INPUT CLAMPS TO RAILS,
* CMRR WITH FREQUENCY EFFECTS, PSRR WITH FREQUENCY EFFECTS,
* SLEW RATE, OPEN LOOP OUTPUT IMPEDANCE, SETTLING TIME TO
* 0.01 PERCENT, QUIESCENT CURRENT WITH TEMPCO, OUTPUT
* CURRENT THROUGH SUPPLIES, OUTPUT CURRENT LIMIT, OUTPUT
* CLAMPS TO RAILS, OUTPUT SWING, OVERLOAD RECOVERY TIME,
* AND OUTPUT OVERSHOOT VERSUS CLOAD
* END MODEL FEATURES
* BEGIN SIMULATION NOTES
* FOR MORE ACCURATE INPUT BIAS CURRENT YOU MAY WANT TO SET
* GMIN FROM THE DEFAULT OF 1E-12 TO 1E-13
* FOR AID IN DC CONVERGENCE SET ITL1 FROM 400 TO 4000
* FOR AID IN TRANSIENT ANALYSIS SET ITL4 FROM 50 TO 500
* MODEL TEMPERATURE RANGE IS -40 C TO +125 C
* NOT ALL PARAMETERS TRACK THOSE OF THE REAL PART VS TEMP
* END SIMULATION NOTES
Q26 8 9 10 QON
Q27 11 9 12 QOP
Q28 13 14 15 QOP 23
Q29 16 17 18 QON 23
I4 8 17 5E-5
I5 14 11 5E-5
R34 19 18 1
R35 15 19 1
R47 20 19 7
E25 11 0 4 0 1
E26 8 0 7 0 1
I9 7 4 3.55E-3
R65 4 7 325E3
R67 12 17 1
R68 14 10 1
R70 21 22 2250
R71 23 22 2250
I11 8 24 5.25E-4
D5 25 8 DD
V9 25 26 -0.4
D6 27 26 DD
V10 27 11 -0.4
E27 28 11 29 11 0.505
C9 9 28 1E-12
R75 28 9 1E3
G2 9 28 30 28 -1E-3
G3 26 28 23 21 -0.19E-3
R76 28 26 1.4E9
C10 30 31 6E-12
R77 30 26 2.2K
E28 32 28 30 28 1
D7 33 34 DD
R78 28 31 220
D8 35 36 DD
C11 21 23 0.4E-12
C12 37 0 4.5E-12
C13 2 0 4.5E-12
L3 20 6 1E-9
R95 6 20 100
E29 32 33 38 0 -2
E30 32 36 38 0 2
R96 33 34 1E12
R97 36 35 1E12
D9 39 0 DD
I12 0 39 1M
R98 38 0 1E12
V11 39 38 0.655
V12 7 16 2.68
V13 13 4 2.68
E42 40 0 41 0 0.023
R113 8 29 1E9
C25 40 29 1E-9
E43 42 0 8 0 0.023
C26 42 41 1E-9
R114 0 41 1E9
E44 43 0 8 0 1
E45 44 0 11 0 1
E46 45 0 46 0 1
R115 43 47 1E6
R116 44 48 1E6
R117 45 49 1E6
R118 0 47 10
R119 0 48 10
R120 0 49 10
E47 50 51 49 0 0.026
R121 52 46 1E3
R122 46 53 1E3
C27 43 47 1E-12
C28 44 48 1E-12
C29 45 49 1E-12
E48 54 50 48 0 -0.06
E49 55 54 47 0 0.01
R123 54 55 1E9
R124 50 54 1E9
R125 51 50 1E9
E50 52 0 2 0 1
E51 53 0 55 0 1
D37 56 57 DL
V145 57 0 3
R316 0 56 1E8
G54 2 0 56 0 2E-10
I67 2 0 5E-12
G55 37 0 56 0 2E-10
I68 37 0 5E-12
D38 58 0 DIN
D39 59 0 DIN
I69 0 58 1E-3
I70 0 59 1E-3
G56 2 55 58 59 2E-11
G57 2 55 60 0 2.4E-7
R317 0 60 1E4
R318 0 60 1E4
D40 61 0 DVN
D41 62 0 DVN
I71 0 61 1E-3
I72 0 62 1E-3
E52 37 55 61 62 0.31
R319 55 37 1E9
V146 26 35 -0.2
V147 34 26 -0.2
V148 63 11 0
V149 8 22 0
J5 64 37 64 JC
J6 64 2 64 JC
V150 8 64 0.25
J7 55 65 55 JC
J8 2 65 2 JC
V151 65 11 0.25
E53 51 66 38 0 5.61E-4
R320 66 51 1E9
V152 66 3 62E-6
G58 7 4 38 0 -6E-3
D42 4 6 DD
D43 6 7 DD
R321 67 68 70
R322 67 69 70
Q30 70 24 63 QIS
Q31 24 24 63 QIS
V153 67 70 0.7
M1 21 37 68 68 NI L=30U W=300U
M2 23 2 69 69 NI L=30U W=300U
M4 71 67 72 72 NS L=30U W=300U
V157 8 73 4.9
R327 71 8 1E5
E55 8 74 8 71 1
R330 73 72 1E3
Q32 9 75 8 QSP
R331 75 74 1E4
C30 55 2 0.45E-12
.MODEL DD D
.MODEL DVN D KF=2.5E-15
.MODEL DIN D KF=1E-15
.MODEL DL D IS=0.95E-11 N=1.4 XTI=1.5
.MODEL NI NMOS VTO=2 KP=1200U IS=1E-18
.MODEL NS NMOS VTO=0 KP=1200U IS=1E-18
.MODEL QSP PNP
.MODEL QIS NPN
.MODEL JC NJF IS=1E-18
.MODEL QON NPN BF=1400 RC=25 TF=150P CJC=100F
.MODEL QOP PNP BF=1400 RC=25 TF=150P CJC=100F
.ENDS OPA827

.param cur=10p
.param offsetv=-0.000071
.param supplyv=15

V_I$3157 POS2 0 offsetv
V_I$1272 POS1 0 offsetv
V_I$1475 VCCP 0 supplyv
V_I$1476 VCCM 0 '-supplyv'
V_I$3150 N$4493 0 supplyv
V_I$3159 N$4492 0 '-supplyv'
L_I$2539 N$2853 N$2855  100p
R_I$2540 N$2855 WE 100
R_I$412 N$2852 N$2853 1k
R_I$208 WE out1 1Meg
R_I$2948 out1 N$4085 0.1K
R_I$3155 N$4085 out2 1Meg
C_I$2542 WE 0 10f
C_I$2541 N$2855 0 10f
C_I$1882 N$2852 N$2853 5f
X_I$5186_I$1 POS2 N$4085 N$4493 N$4492 out2  OPA827 
X_I$4984_I$1 POS1 WE VCCP VCCM out1  OPA827 
I_I$411 0 N$2852 pwl(0 0 1 100p)

.trans 1u 1
.extract label=vmax1 max(v(out1))
.extract label=vmin1 min(v(out1))
.extract label=vmax2 max(v(out2))
.extract label=vmin2 min(v(out2))
.plot v(out1)
.plot v(out2)
.plot i(I_I$411)

.op  NO_SMALL_SIGNAL
.END
